* EBeam Silicon photonic circuit
*
  
.subckt Simple_MZI N$0 N$1
	Xebeam_gc_te1550_0 N$0 N$2 ebeam_gc_te1550 library="Design kits/ebeam_v1.0" sch_x=150.0e-3 sch_y=700.0e-3 
	Xebeam_gc_te1550_1 N$1 N$3 ebeam_gc_te1550 library="Design kits/ebeam_v1.0" sch_x=150.0e-3 sch_y=7.05 
	Xebeam_y_1550_2 N$4 N$5 N$6 ebeam_y_1550 library="Design kits/ebeam_v1.0" sch_x=2.0 sch_y=6.2 
	Xebeam_y_1550_3 N$7 N$8 N$9 ebeam_y_1550 library="Design kits/ebeam_v1.0" sch_x=2.0 sch_y=1.45 
	Xwg0 N$3 N$4 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" wg_length=54.1e-6 wg_width=500.0e-9 	sch_x=1.11625 sch_y=6.625
	Xwg1 N$6 N$8 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" wg_length=133.5e-6 wg_width=500.0e-9 	sch_x=3.3 sch_y=3.825
	Xwg2 N$9 N$5 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" wg_length=154.5e-6 wg_width=500.0e-9 	sch_x=3.425 sch_y=3.825
	Xwg3 N$7 N$2 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" wg_length=52.1e-6 wg_width=500.0e-9 	sch_x=916.25e-3 sch_y=1.075
.ends Simple_MZI

* - ONA
.ona input_unit=wavelength input_parameter=center_and_range center=1550e-9
  + range=100e-9 number_of_points=3000 
  + minimum_loss=50
  + sensitivity=-200 
  + analysis_type=scattering_data
  + multithreading=user_defined number_of_threads=1 
  + input(1)=Simple_MZI,N$0
  + output=Simple_MZI,N$1

Simple_MZI N$0 N$1 Simple_MZI sch_x=-1 sch_y=-1

.end
