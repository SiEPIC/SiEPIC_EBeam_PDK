* Spice output from KLayout SiEPIC_EBeam_PDK v0.1.6, 2015-11-26 01:30:46.

.subckt wg_test2
  x0  N$0 "Waveguide Arc Bend" library="Waveguides/Bends" lay_x=-53.0u lay_y=21.4u sch_x=-10.6 sch_y=4.28  sch_r=450 sch_f=true
  x1  N$1 N$2 "Waveguide Arc Bend" library="Waveguides/Bends" lay_x=10.8u lay_y=21.4u sch_x=2.16 sch_y=4.28  sch_r=360 sch_f=true
  x2  N$3 N$4 "Waveguide Arc Bend" library="Waveguides/Bends" lay_x=10.8u lay_y=-67.0u sch_x=2.16 sch_y=-13.4  sch_r=270
  x3  N$5 N$6 "Waveguide Arc Bend" library="Waveguides/Bends" lay_x=74.2u lay_y=-67.0u sch_x=14.84 sch_y=-13.4 
  x4  N$7 N$8 "Waveguide Arc Bend" library="Waveguides/Bends" lay_x=74.2u lay_y=20.2u sch_x=14.84 sch_y=4.04  sch_r=450 sch_f=true
  x5  N$9 "Waveguide Arc Bend" library="Waveguides/Bends" lay_x=152.9u lay_y=20.2u sch_x=30.58 sch_y=4.04  sch_r=360 sch_f=true
  x6  N$0 N$1 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" lay_x=-21.1u lay_y=21.4u sch_x=-4.22 sch_y=4.28 
  x7  N$2 N$3 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" lay_x=10.8u lay_y=-22.8u sch_x=2.16 sch_y=-4.56  sch_r=270
  x8  N$4 N$5 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" lay_x=42.5u lay_y=-67.0u sch_x=8.5 sch_y=-13.4 
  x9  N$6 N$7 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" lay_x=74.2u lay_y=-23.4u sch_x=14.84 sch_y=-4.68  sch_r=90
  x10  N$8 N$9 ebeam_wg_strip_1550 library="Design kits/ebeam_v1.0" lay_x=113.55u lay_y=20.2u sch_x=22.71 sch_y=4.04 
.ends wg_test2

wg_test2 wg_test2 sch_x=-1 sch_y=-1

